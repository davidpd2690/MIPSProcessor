module ForwardingUnit
(
	input IDEX_RegisterRs,
	input IDEX_RegisterRt,
	
	input EXMEM_RegWrite,
	input EXMEM_RegisterRd,
	
	input MEMWB_RegWrite,
	input MEMWB_RegisterRd,
	
	output ForwardA,
	output ForwardB
);





endmodule